`ifndef __TEST_TOP_SV_
`define __TEST_TOP_SV_

`include "base_test.sv"

`include "random_data_add_test.sv"
`include "order_data_add_test.sv"
`include "burst_nodelay_add_test.sv"
`include "random_delay_add_test.sv"

`endif
